// ============================================================
// Q1.15 Trig LUT ROM for Hough Transform
// - Loads sine/cosine tables from .mem files
// - Inferred as M9K BRAMs (DE2 Cyclone II)
// ============================================================
module trig_lut_rom #(
    parameter THETA_STEPS = 180
)(
    input  logic clk,
    input  logic [$clog2(THETA_STEPS)-1:0] theta_idx,
    output logic signed [15:0] cos_q,
    output logic signed [15:0] sin_q
);

    // ------------------------------------------------------------
    // M9K block RAM inference
    // ------------------------------------------------------------
    (* ramstyle = "M9K", romstyle = "M9K" *) reg signed [15:0] cos_rom [0:THETA_STEPS-1];
    (* ramstyle = "M9K", romstyle = "M9K" *) reg signed [15:0] sin_rom [0:THETA_STEPS-1];

    // ------------------------------------------------------------
    // Load data from external .mem files (generated by Python)
    // ------------------------------------------------------------
    initial begin
        $readmemh("cos_lut.mem", cos_rom);
        $readmemh("sin_lut.mem", sin_rom);
    end

    // ------------------------------------------------------------
    // 1-cycle latency synchronous read
    // ------------------------------------------------------------
    always_ff @(posedge clk) begin
        cos_q <= cos_rom[theta_idx];
        sin_q <= sin_rom[theta_idx];
    end

endmodule
// ============================================================
