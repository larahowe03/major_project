// hi tumali